module acceleratorTB;


endmodule
